module decoder1();
